��u       �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�base_estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.0.1�ub�n_estimators�K
�estimator_params�(hhhhhhhhhht��	bootstrap���	oob_score���n_jobs�NhK �verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        h�auto�hNhG        hG        �feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h)�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�objawy��wiek��choroby��wzrost�et�b�n_features_in_�K�
n_outputs_�K�classes_�h(h+K ��h-��R�(KK��h2�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�base_estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hh$hNhJ�
hG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��h2�f8�����R�(KhHNNNJ����J����K t�b�C              �?�t�bhLh&�scalar���hGC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hK�
node_count�K�nodes�h(h+K ��h-��R�(KK��h2�V56�����R�(Kh6N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hxhGK ��hyhGK��hzhGK��h{hXK��h|hXK ��h}hGK(��h~hXK0��uK8KKt�b�B                              @*O���?             B@                           @ �q�q�?             8@������������������������       �                     7@������������������������       �                     �?������������������������       �        
             (@�t�b�values�h(h+K ��h-��R�(KKKK��hX�CP      7@      *@      7@      �?      7@                      �?              (@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ/��hG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoKhph(h+K ��h-��R�(KK��hw�C�                            @X�<ݚ�?             B@������������������������       �                     0@������������������������       �                     4@�t�bh�h(h+K ��h-��R�(KKKK��hX�C0      0@      4@      0@                      4@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJu�7hG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoKhph(h+K ��h-��R�(KK��hw�B�                              @)O���?             B@������������������������       �                     1@                            @�KM�]�?             3@                           @���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     ,@�t�bh�h(h+K ��h-��R�(KKKK��hX�Cp      3@      1@      1@               @      1@       @      @       @                      @              ,@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��!XhG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoKhph(h+K ��h-��R�(KK��hw�B�                              @X�<ݚ�?             B@                           P@�C��2(�?             6@������������������������       �                     3@                            @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     ,@�t�bh�h(h+K ��h-��R�(KKKK��hX�Cp      4@      0@      4@       @      3@              �?       @      �?                       @              ,@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJC�NhG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoKhph(h+K ��h-��R�(KK��hw�B�                              @�q�q�?             B@                            @���7�?             6@������������������������       �                     2@                         yJK@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     ,@�t�bh�h(h+K ��h-��R�(KKKK��hX�Cp      5@      .@      5@      �?      2@              @      �?      @                      �?              ,@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�R�[hG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoKhph(h+K ��h-��R�(KK��hw�B�                           �%g@X�<ݚ�?             B@                           @ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?                            @
j*D>�?             :@������������������������       �                     &@������������������������       �                     .@�t�bh�h(h+K ��h-��R�(KKKK��hX�Cp      4@      0@      "@      �?      "@                      �?      &@      .@      &@                      .@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�v}hG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoKhph(h+K ��h-��R�(KK��hw�B�                            pg@)O���?             B@                            @d}h���?	             ,@������������������������       �                     &@������������������������       �                     @                            @���!pc�?             6@������������������������       �                     @������������������������       �                     0@�t�bh�h(h+K ��h-��R�(KKKK��hX�Cp      1@      3@      &@      @      &@                      @      @      0@      @                      0@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJg}�XhG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoKhph(h+K ��h-��R�(KK��hw�B                              @      �?             B@                           @؇���X�?             5@������������������������       �                     2@������������������������       �                     @������������������������       �        
             .@�t�bh�h(h+K ��h-��R�(KKKK��hX�CP      2@      2@      2@      @      2@                      @              .@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ	�tlhG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoKhph(h+K ��h-��R�(KK��hw�B                            �e@)O���?             B@������������������������       �                     @                            @J�8���?             =@������������������������       �                     $@������������������������       �                     3@�t�bh�h(h+K ��h-��R�(KKKK��hX�CP      1@      3@      @              $@      3@      $@                      3@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�ޡhG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoKhph(h+K ��h-��R�(KK��hw�C�                            @)O���?             B@������������������������       �                     3@������������������������       �                     1@�t�bh�h(h+K ��h-��R�(KKKK��hX�C0      3@      1@      3@                      1@�t�bubhhubehhub.